* Analog to Manchester Encoder
* Design by: Skull0nFire
* Wed, Apr 28, 2021 02:22:43 
********************
*INPUTS FOR TESTING*
********************
vin     inp 0 sine(2    2   50  0   0   0)
vSL     SL  0 PULSE(0   5   2m  1n  1n  2.66m   4m)
vclk    clk 0 PULSE(0   5   0   1n  1n  0.66m   1.33m)

.include ua741.cir
.include ADC8bit.cir
.include PISO.cir

*******************************
*Manchester Encoder Subcircuit*
*******************************
.subckt ManchesterEnc   inp SL  clk sout manchester 
*****************************************************************************
*Connecting the ADC, PISO and XOR gate to get the required Manchester Signal*
*****************************************************************************
Xu1 inp out0    out1    out2    v1  v2  v3  v4  v5  v6  v7  ADC8bit

Xu2 SL  clk     out0    out1    out2    sout    PISO

Xu3 clk sout    manchester  xor
.ends   ManchesterEnc


Xu0 inp SL  clk sout    manchester  ManchesterEnc

.tran 10u 50m
.control
run

set color0=white
set color1=black 
set color2=red
set color3=darkorange
set color4=Teal
set color5=darkblue
set color6=darkgreen
set color7=magenta
set Xbrushwidth=2

plot    v(inp)
plot    v(clk)  v(SL)+5.5   v(sout)+11  v(manchester)+16.5

.endc
.end