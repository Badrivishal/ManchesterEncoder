*Parallel IN Serial OUT
********************
*INPUTS FOR TESTING*
********************
* vb0 b0 0 PULSE(0 5 1m 0 0 4m 8m)
* vb1 b1 0 PULSE(0 5 1m 0 0 8m 16m)
* vb2 b2 0 PULSE(0 5 1m 0 0 16m 32m)
* vSL SL 0 PULSE(0 5 2m 0 0 2.66m 4m)
* vclk clk 0 PULSE(0 5 0 0 0 0.66m 1.33m)

.include AOI_BasicGatesCkts.cir

****************
*3 inp NOR gate*
****************
.subckt nor3 in1 in2 in3 out
Xn1 in1 in2 n0 nor
Xn2 n0 n0 n1 nor
Xn3 n1 in3 out nor
.ends


************************************
*Negative edge triggered D flipFlop*
************************************
.subckt flipFlopD d clk q notq

X4 n0 d n1 nor
X3 n3 clk n1 n0 nor3
X2 n2 clk n3 nor
X1 n1 n3 n2 nor

X5 n3 notq q nor
X6 q n0 notq nor
.ends

***********************
*3 BIT PISO SUBCIRCUIT*
***********************
.subckt PISO SL clk b0 b1 b2 q2
Xn1 SL notSL not

Xd0 b0 clk q0 notq0 flipFlopD

Xa1 q0 SL n0 and
Xa2 notSL b1 n1 and
Xo1 n0 n1 d1 or

Xd1 d1 clk q1 notq1 flipFlopD

Xa3 q1 SL n2 and
Xa4 notSL b2 n3 and
Xo2 n2 n3 d2 or

Xd2 d2 clk q2 notq2 flipFlopD

.ends PISO


* Xu1 SL clk b0 b1 b2 q2 PISO

* .tran 10u 32m 
* .control
* run

* set color0=black
* set color1=white
* set color2=red
* set color3=blue
* set color4=green
* set Xbrushwidth=2

* plot v(clk) v(SL)+5 v(q2)+10
* plot v(b0) v(b1) v(b2)
.endc
.end
